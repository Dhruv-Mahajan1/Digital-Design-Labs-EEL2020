`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/04/2022 07:13:41 PM
// Design Name: 
// Module Name: TestCarryLookAhead
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TestCarryLookAhead();
reg [31:0] A,B;
reg Cin;
wire [31:0]OutputSum;
wire Cout;
CarryLookAhead CLA(A,B,Cin,OutputSum,Cout);
initial
    begin
        Cin=1'b0;
        A=32'b00000000000000000000000000000000; B=32'b00000000000000000000000000000000;
        #10 A=32'b00000000000000000000000000000010; B=32'b00000000000000000000000000000001;
        #10 A=32'b00000000000000000000000000001000; B=32'b00000000000000000000000000000010;
        #10 A=32'b00000000000000000000000000100000; B=32'b00000000000000000000000100000000;
        #10 A=32'b00000000000000000000000000000000; B=32'b00000000000000000000000000000000;
        #10 A=32'b00000000000000000001000000000000; B=32'b00000000000000000000000001000000;
        #10 A=32'b00000000000000000000000001000000; B=32'b00000000001000000000000000000000;
        #10 A=32'b00000000000000000100000000000000; B=32'b00000001000000000000000000000000;
        #10 A=32'b00000000000000000001000000000000; B=32'b00000000000000000000000000100000;
        #10 A=32'b00000000000010000000000000000000; B=32'b00000000001000000000000000000000;
        #10 A=32'b00000000000000000000000001000000; B=32'b00000000000000000000000010000000;
       
        
    end

initial #110 $finish;
endmodule

